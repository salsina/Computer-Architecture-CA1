module tb();
    reg [5:0] x,y;
    wire [11:0] result;
    reg clk,rst,start;
    wire ldx,ldy,shiftY,init_result,initcnt,encnt,ldresult,en_mult_one_bit_y,carryout;
    wire done;
    datapath dp(x,y,ldx,ldy,shiftY,clk,rst,initcnt,encnt,en_mult_one_bit_y,init_result,ldresult,result,carryout);
    controller cntlr(clk,rst,carryout,start,ldx,ldy,shiftY,initcnt,encnt,en_mult_one_bit_y,init_result,ldresult,done);
initial begin
        start=0; x=-16; y=5; rst=1;
        clk=0;
        #20 clk=1;
        #20 clk=0; rst=0;
        start=1;
        #20 clk=0;
        #20 clk=1;
        #20 clk=0;
        #20 clk=1;
        #20 clk=0;
        start = 0;
        #20 clk=1;
        #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
        #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
        #20 clk=0;
        x=-25; y=-4;
        #20 clk=1;
        #20 clk=0; rst=0;
        start=1;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        start = 0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
        #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
	    #20 clk=0;
        #20 clk=1;
        #200;
    end
endmodule